/*
	a simple program to demonstrate the use of and gate
*/
module combin (
	input in1,
	input in2,
	output out
	);

	assign out = in1 & in2;

endmodule
